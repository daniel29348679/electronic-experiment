`timescale 1ns / 1ps
module TM;

    reg clk;

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    reg reset;
    wire [3:0] count;

    Counter counter (
        .clk (clk),
        .rst (reset),
        .dout(count)
    );

    integer i;

    initial begin
        $dumpfile("test.vcd");
        $dumpvars(0, counter);
        $monitor("reset = %b, count = %d", reset, count);
        for (i = 0; i < 200; i = i + 1) begin
            reset <= (i % 11 == 0);
            #10;
        end
        $finish;

    end
endmodule
